
module lc_ulpb_bridge(DATA_FROM_LC, ADDR_FROM_LC, REQ_FROM_LC, ACK_TO_LC,
					  DATA_TO_LC, ADDR_TO_LC, REQ_TO_LC, ACK_FROM_LC,
					  CLK, RESET, REQ_TX, DATA_BUF1, DATA_BUF2, DATA_PENDING, ADDR_OUT, DATA_INDICATOR)

input	CLK, RESET;

parameter DATA_WIDTH=32;
parameter ADDR_WIDTH=8;

input	[ADDR_WIDTH-1:0] ADDR_FROM_LC;
input	[DATA_WIDTH-1:0] DATA_FROM_LC;
input	REQ_FROM_LC;
output	ACK_TO_LC;

output  [ADDR_WIDTH-1:0] ADDR_TO_LC;
output  [DATA_WIDTH-1:0] DATA_TO_LC;
output  REQ_TO_LC;
input	ACK_FROM_LC;

output	REQ_TX;
output	[DATA_WIDTH-1:0] DATA_BUF1, DATA_BUF2;
output	[ADDR_WIDTH-1:0] ADDR_OUT;
output	DATA_PENDING;
input	DATA_INDICATOR;
