// Verilog HDL and netlist files of
// "SLEEP_CONTROL SLEEP_CONTROLv4 schematic"

// Library - SLEEP_CONTROL, Cell - SLEEP_CONTROLv4, View - schematic
// LAST TIME SAVED: Apr 10 15:16:23 2013
// NETLIST TIME: Apr 10 15:41:53 2013
`timescale 1ns / 1ns 
`include "/afs/eecs.umich.edu/kits/ARM/TSMC_cl018g/mosis_2009q1/sc-x_2004q3v1/aci/sc/verilog/tsmc18_neg.v"

module SLEEP_CONTROLv4 ( MBC_ISOLATE, MBC_ISOLATE_B, MBC_RESET,
     MBC_RESET_B, MBC_SLEEP, MBC_SLEEP_B, SYSTEM_ACTIVE,
     WAKEUP_REQ_ORED, /*VDD, VSS,*/ CLK, MBUS_DIN, RESETn, SLEEP_REQ,
     WAKEUP_REQ0, WAKEUP_REQ1, WAKEUP_REQ2 );

output  MBC_ISOLATE, MBC_ISOLATE_B, MBC_RESET, MBC_RESET_B, MBC_SLEEP,
     MBC_SLEEP_B, SYSTEM_ACTIVE, WAKEUP_REQ_ORED;

//inout  VDD, VSS;

input  CLK, MBUS_DIN, RESETn, SLEEP_REQ, WAKEUP_REQ0, WAKEUP_REQ1,
     WAKEUP_REQ2;


NOR3X1 I1 ( .C(WAKEUP_REQ2), .B(WAKEUP_REQ1), .A(WAKEUP_REQ0), .Y(WAKEUP_REQ_ORED_B_int) );
INVX2 I2 ( .Y(WAKEUP_REQ_ORED), .A(WAKEUP_REQ_ORED_B_int));
INVX1 I27 ( .Y(net071), .A(net02));
INVX1 I13 ( .Y(RESET), .A(RESETn));
INVX1 I10 ( .Y(MBUS_DIN_B), .A(MBUS_DIN));
INVX1 I3 ( .Y(SLEEP_REQ_B), .A(SLEEP_REQ));
DFFSRX1 I19 ( .SN(RESETn), .RN(VDD), .CK(CLK), .Q(MBC_RESET_int), .QN(MBC_RESET_B_int), .D(MBC_ISOLATE_int));
DFFSRX1 I15 ( .SN(RESETn), .RN(VDD), .CK(CLK), .Q(MBC_ISOLATE_int), .QN(MBC_ISOLATE_B_int), .D(net057));
DFFSRX1 I7 ( .SN(SETn_TRAN_TO_WAKE), .RN(RSTn_TRAN_TO_WAKE), .CK(VSS),   .Q(TRAN_TO_WAKE), .QN(net035), .D(VSS));
DFFSRX1 I4 ( .SN(RESETn), .RN(VDD), .CK(CLK), .Q(MBC_SLEEP_int), .QN(MBC_SLEEP_B_int), .D(net014));
NAND2X1 I29 ( .Y(SYSTEM_ACTIVE), .A(MBC_SLEEP), .B(MBC_ISOLATE_int));
NAND2X1 I22 ( .Y(net057), .A(TRAN_TO_WAKE), .B(MBC_SLEEP_B_int));
NAND2X1 I11 ( .Y(net034), .A(MBC_SLEEP_int), .B(MBUS_DIN_B));
NAND2X1 I9 ( .Y(SET_TRAN_TO_WAKE_ifnoporeset), .A(WAKEUP_REQ_ORED_B_int), .B(net034));
NAND2X1 I8 ( .B(RESETn), .A(SET_TRAN_TO_WAKE_ifnoporeset), .Y(SETn_TRAN_TO_WAKE), .VSS(VSS));
NOR2X1 I26 ( .B(MBC_SLEEP_B_int), .A(SET_TRAN_TO_WAKE_ifnoporeset), .Y(net02), .VSS(VSS));
NOR2X1 I21 ( .B(MBC_ISOLATE_B_int), .A(TRAN_TO_WAKE), .Y(net014), .VSS(VSS));
NOR2X1 I14 ( .B(SLEEP_REQ_B), .A(SET_TRAN_TO_WAKE_ifnoporeset), .Y(net033), .VSS(VSS));
NOR2X1 I12 ( .Y(RSTn_TRAN_TO_WAKE), .A(net033), .B(RESET));
INVX12 I28 ( .Y(MBC_SLEEP_B), .A(net02));
INVX12 I25 ( .Y(MBC_ISOLATE_B), .A(MBC_ISOLATE_int));
INVX12 I24 ( .Y(MBC_RESET_B), .A(MBC_RESET_int));
INVX12 I23 ( .Y(MBC_SLEEP), .A(net071));
INVX12 I20 ( .Y(MBC_RESET), .A(MBC_RESET_B_int));
INVX12 I18 ( .Y(MBC_ISOLATE), .A(MBC_ISOLATE_B_int));

endmodule


// End HDL models
